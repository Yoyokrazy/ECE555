* SPICE NETLIST
***************************************

.SUBCKT NEURON VSS VDD X_1<0> X_0<0> W1_0<0> W1_0<1> W0_0<0> W0_0<1> X_1<1> X_0<1> CIN_0 W2_0<0> W2_0<1> W2_0<2> CIN_1 COUT Z<2> Z<1> Z<0>
** N=430 EP=19 IP=0 FDC=298
M0 11 X_1<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=972 $D=0
M1 VDD 4 15 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=1512 $D=0
M2 12 X_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=3456 $D=0
M3 VDD 6 16 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=3996 $D=0
M4 VDD W1_0<0> 11 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=972 $D=0
M5 142 W1_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=1512 $D=0
M6 VDD W0_0<0> 12 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=3456 $D=0
M7 143 W0_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=3996 $D=0
M8 15 X_1<1> 142 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=1512 $D=0
M9 16 X_0<1> 143 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=3996 $D=0
M10 19 11 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1296 $Y=972 $D=0
M11 20 12 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1296 $Y=3456 $D=0
M12 4 X_1<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=1512 $D=0
M13 6 X_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=3996 $D=0
M14 VDD W1_0<1> 4 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=1512 $D=0
M15 VDD W0_0<1> 6 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=3996 $D=0
M16 17 15 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=1512 $D=0
M17 18 16 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=3996 $D=0
M18 21 17 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=972 $D=0
M19 VDD 15 17 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=1512 $D=0
M20 22 18 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=3456 $D=0
M21 VDD 16 18 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=3996 $D=0
M22 VDD 19 21 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=972 $D=0
M23 VDD 20 22 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=3456 $D=0
M24 24 21 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3024 $Y=972 $D=0
M25 26 22 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3024 $Y=3456 $D=0
M26 27 20 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=972 $D=0
M27 VDD 23 29 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=1512 $D=0
M28 28 24 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=3456 $D=0
M29 VDD 25 30 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=3996 $D=0
M30 VDD 19 27 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=972 $D=0
M31 144 20 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=1512 $D=0
M32 VDD 26 28 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=3456 $D=0
M33 145 24 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=3996 $D=0
M34 29 19 144 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=1512 $D=0
M35 30 26 145 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=3996 $D=0
M36 41 27 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4752 $Y=972 $D=0
M37 42 28 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4752 $Y=3456 $D=0
M38 23 19 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=1512 $D=0
M39 25 26 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=3996 $D=0
M40 VDD 20 23 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=1512 $D=0
M41 VDD 24 25 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=3996 $D=0
M42 31 29 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=1512 $D=0
M43 32 30 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=3996 $D=0
M44 37 31 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5616 $Y=972 $D=0
M45 VDD 29 31 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=1512 $D=0
M46 38 32 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5616 $Y=3456 $D=0
M47 VDD 30 32 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=3996 $D=0
M48 VDD CIN_0 37 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5832 $Y=972 $D=0
M49 VDD 34 38 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5832 $Y=3456 $D=0
M50 VDD 35 43 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=1512 $D=0
M51 VDD 36 44 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=3996 $D=0
M52 39 37 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6480 $Y=972 $D=0
M53 146 CIN_0 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=1512 $D=0
M54 40 38 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6480 $Y=3456 $D=0
M55 147 34 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=3996 $D=0
M56 43 31 146 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=1512 $D=0
M57 44 32 147 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=3996 $D=0
M58 117 39 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7128 $Y=972 $D=0
M59 118 40 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7128 $Y=3456 $D=0
M60 45 41 117 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=972 $D=0
M61 35 31 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=1512 $D=0
M62 46 42 118 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=3456 $D=0
M63 36 32 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=3996 $D=0
M64 VDD CIN_0 35 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7560 $Y=1512 $D=0
M65 VDD 34 36 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7560 $Y=3996 $D=0
M66 53 43 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=1512 $D=0
M67 54 44 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=3996 $D=0
M68 34 45 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7992 $Y=972 $D=0
M69 VDD 43 53 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=1512 $D=0
M70 55 46 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7992 $Y=3456 $D=0
M71 VDD 44 54 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=3996 $D=0
M72 56 W2_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=972 $D=0
M73 VDD 48 59 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=1512 $D=0
M74 57 W2_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=3456 $D=0
M75 VDD 50 60 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=3996 $D=0
M76 58 W2_0<2> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=5940 $D=0
M77 VDD 52 61 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=6480 $D=0
M78 VDD 53 56 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=972 $D=0
M79 148 W2_0<0> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=1512 $D=0
M80 VDD 54 57 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=3456 $D=0
M81 149 W2_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=3996 $D=0
M82 VDD 55 58 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=5940 $D=0
M83 150 W2_0<2> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=6480 $D=0
M84 59 53 148 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=1512 $D=0
M85 60 54 149 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=3996 $D=0
M86 61 55 150 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=6480 $D=0
M87 77 56 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10016 $Y=972 $D=0
M88 78 57 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10016 $Y=3456 $D=0
M89 79 58 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10016 $Y=5940 $D=0
M90 48 53 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=1512 $D=0
M91 50 54 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=3996 $D=0
M92 52 55 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=6480 $D=0
M93 VDD W2_0<0> 48 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=1512 $D=0
M94 VDD W2_0<1> 50 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=3996 $D=0
M95 VDD W2_0<2> 52 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=6480 $D=0
M96 62 59 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=1512 $D=0
M97 63 60 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=3996 $D=0
M98 64 61 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=6480 $D=0
M99 71 62 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=972 $D=0
M100 VDD 59 62 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=1512 $D=0
M101 72 63 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=3456 $D=0
M102 VDD 60 63 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=3996 $D=0
M103 73 64 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=5940 $D=0
M104 VDD 61 64 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=6480 $D=0
M105 VDD CIN_1 71 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=972 $D=0
M106 VDD 66 72 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=3456 $D=0
M107 VDD 67 73 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=5940 $D=0
M108 VDD 68 80 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=1512 $D=0
M109 VDD 69 81 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=3996 $D=0
M110 VDD 70 82 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=6480 $D=0
M111 74 71 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11744 $Y=972 $D=0
M112 151 CIN_1 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=1512 $D=0
M113 75 72 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11744 $Y=3456 $D=0
M114 152 66 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=3996 $D=0
M115 76 73 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11744 $Y=5940 $D=0
M116 153 67 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=6480 $D=0
M117 80 62 151 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=1512 $D=0
M118 81 63 152 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=3996 $D=0
M119 82 64 153 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=6480 $D=0
M120 125 74 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=972 $D=0
M121 126 75 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=3456 $D=0
M122 127 76 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=5940 $D=0
M123 83 77 125 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=972 $D=0
M124 68 62 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=1512 $D=0
M125 84 78 126 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=3456 $D=0
M126 69 63 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=3996 $D=0
M127 85 79 127 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=5940 $D=0
M128 70 64 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=6480 $D=0
M129 VDD CIN_1 68 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=1512 $D=0
M130 VDD 66 69 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=3996 $D=0
M131 VDD 67 70 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=6480 $D=0
M132 89 80 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=1512 $D=0
M133 88 81 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=3996 $D=0
M134 86 82 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=6480 $D=0
M135 66 83 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=972 $D=0
M136 VDD 80 89 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=1512 $D=0
M137 67 84 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=3456 $D=0
M138 VDD 81 88 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=3996 $D=0
M139 COUT 85 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=5940 $D=0
M140 VDD 82 86 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=6480 $D=0
M141 Z<2> VDD VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=14464 $Y=3696 $D=0
M142 87 86 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=14464 $Y=4236 $D=0
M143 90 87 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=15408 $Y=3804 $D=0
M144 91 88 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=15408 $Y=4236 $D=0
M145 VDD 89 90 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=15624 $Y=3804 $D=0
M146 VDD 87 91 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=15624 $Y=4236 $D=0
M147 Z<1> 90 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=16272 $Y=3804 $D=0
M148 Z<0> 91 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=16272 $Y=4236 $D=0
M149 109 X_1<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=108 $D=1
M150 92 4 15 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=2052 $D=1
M151 110 X_0<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=2592 $D=1
M152 93 6 16 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=4536 $D=1
M153 11 W1_0<0> 109 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=108 $D=1
M154 VSS W1_0<1> 92 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=2052 $D=1
M155 12 W0_0<0> 110 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=2592 $D=1
M156 VSS W0_0<1> 93 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=4536 $D=1
M157 92 X_1<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=2052 $D=1
M158 93 X_0<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=4536 $D=1
M159 19 11 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=108 $D=1
M160 20 12 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=2592 $D=1
M161 130 X_1<1> 4 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=2052 $D=1
M162 131 X_0<1> 6 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=4536 $D=1
M163 VSS W1_0<1> 130 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=2052 $D=1
M164 VSS W0_0<1> 131 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=4536 $D=1
M165 17 15 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=2052 $D=1
M166 18 16 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=4536 $D=1
M167 111 17 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=108 $D=1
M168 VSS 15 17 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=2052 $D=1
M169 112 18 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=2592 $D=1
M170 VSS 16 18 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=4536 $D=1
M171 21 19 111 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=108 $D=1
M172 22 20 112 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=2592 $D=1
M173 24 21 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=108 $D=1
M174 26 22 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=2592 $D=1
M175 113 20 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=108 $D=1
M176 94 23 29 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=2052 $D=1
M177 114 24 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=2592 $D=1
M178 95 25 30 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=4536 $D=1
M179 27 19 113 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4104 $Y=108 $D=1
M180 VSS 20 94 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=2052 $D=1
M181 28 26 114 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4104 $Y=2592 $D=1
M182 VSS 24 95 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=4536 $D=1
M183 94 19 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=2052 $D=1
M184 95 26 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=4536 $D=1
M185 41 27 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=108 $D=1
M186 42 28 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=2592 $D=1
M187 132 19 23 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4968 $Y=2052 $D=1
M188 133 26 25 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4968 $Y=4536 $D=1
M189 VSS 20 132 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5184 $Y=2052 $D=1
M190 VSS 24 133 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5184 $Y=4536 $D=1
M191 31 29 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=2052 $D=1
M192 32 30 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=4536 $D=1
M193 115 31 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5616 $Y=108 $D=1
M194 VSS 29 31 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=2052 $D=1
M195 116 32 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5616 $Y=2592 $D=1
M196 VSS 30 32 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=4536 $D=1
M197 37 CIN_0 115 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5832 $Y=108 $D=1
M198 38 34 116 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5832 $Y=2592 $D=1
M199 96 35 43 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=2052 $D=1
M200 97 36 44 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=4536 $D=1
M201 39 37 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=108 $D=1
M202 VSS CIN_0 96 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=2052 $D=1
M203 40 38 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=2592 $D=1
M204 VSS 34 97 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=4536 $D=1
M205 96 31 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=2052 $D=1
M206 97 32 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=4536 $D=1
M207 45 39 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7128 $Y=108 $D=1
M208 46 40 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7128 $Y=2592 $D=1
M209 VSS 41 45 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7344 $Y=108 $D=1
M210 134 31 35 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7344 $Y=2052 $D=1
M211 VSS 42 46 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7344 $Y=2592 $D=1
M212 135 32 36 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7344 $Y=4536 $D=1
M213 VSS CIN_0 134 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7560 $Y=2052 $D=1
M214 VSS 34 135 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7560 $Y=4536 $D=1
M215 53 43 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=2052 $D=1
M216 54 44 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=4536 $D=1
M217 34 45 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7992 $Y=108 $D=1
M218 VSS 43 53 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=2052 $D=1
M219 55 46 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7992 $Y=2592 $D=1
M220 VSS 44 54 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=4536 $D=1
M221 119 W2_0<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=108 $D=1
M222 99 48 59 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=2052 $D=1
M223 120 W2_0<1> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=2592 $D=1
M224 100 50 60 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=4536 $D=1
M225 121 W2_0<2> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=5076 $D=1
M226 101 52 61 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=7020 $D=1
M227 56 53 119 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=108 $D=1
M228 VSS W2_0<0> 99 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=2052 $D=1
M229 57 54 120 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=2592 $D=1
M230 VSS W2_0<1> 100 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=4536 $D=1
M231 58 55 121 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=5076 $D=1
M232 VSS W2_0<2> 101 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=7020 $D=1
M233 99 53 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=2052 $D=1
M234 100 54 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=4536 $D=1
M235 101 55 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=7020 $D=1
M236 77 56 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=108 $D=1
M237 78 57 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=2592 $D=1
M238 79 58 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=5076 $D=1
M239 136 53 48 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=2052 $D=1
M240 137 54 50 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=4536 $D=1
M241 138 55 52 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=7020 $D=1
M242 VSS W2_0<0> 136 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=2052 $D=1
M243 VSS W2_0<1> 137 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=4536 $D=1
M244 VSS W2_0<2> 138 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=7020 $D=1
M245 62 59 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=2052 $D=1
M246 63 60 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=4536 $D=1
M247 64 61 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=7020 $D=1
M248 122 62 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=108 $D=1
M249 VSS 59 62 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=2052 $D=1
M250 123 63 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=2592 $D=1
M251 VSS 60 63 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=4536 $D=1
M252 124 64 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=5076 $D=1
M253 VSS 61 64 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=7020 $D=1
M254 71 CIN_1 122 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=108 $D=1
M255 72 66 123 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=2592 $D=1
M256 73 67 124 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=5076 $D=1
M257 102 68 80 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=2052 $D=1
M258 103 69 81 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=4536 $D=1
M259 104 70 82 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=7020 $D=1
M260 74 71 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=108 $D=1
M261 VSS CIN_1 102 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=2052 $D=1
M262 75 72 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=2592 $D=1
M263 VSS 66 103 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=4536 $D=1
M264 76 73 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=5076 $D=1
M265 VSS 67 104 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=7020 $D=1
M266 102 62 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=2052 $D=1
M267 103 63 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=4536 $D=1
M268 104 64 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=7020 $D=1
M269 83 74 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=108 $D=1
M270 84 75 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=2592 $D=1
M271 85 76 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=5076 $D=1
M272 VSS 77 83 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=108 $D=1
M273 139 62 68 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=2052 $D=1
M274 VSS 78 84 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=2592 $D=1
M275 140 63 69 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=4536 $D=1
M276 VSS 79 85 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=5076 $D=1
M277 141 64 70 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=7020 $D=1
M278 VSS CIN_1 139 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=2052 $D=1
M279 VSS 66 140 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=4536 $D=1
M280 VSS 67 141 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=7020 $D=1
M281 89 80 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=2052 $D=1
M282 88 81 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=4536 $D=1
M283 86 82 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=7020 $D=1
M284 66 83 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=108 $D=1
M285 VSS 80 89 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=2052 $D=1
M286 67 84 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=2592 $D=1
M287 VSS 81 88 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=4536 $D=1
M288 COUT 85 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=5076 $D=1
M289 VSS 82 86 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=7020 $D=1
M290 Z<2> VDD VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=14464 $Y=2940 $D=1
M291 87 86 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=14464 $Y=4992 $D=1
M292 128 87 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=15408 $Y=2940 $D=1
M293 129 88 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=15408 $Y=4884 $D=1
M294 90 89 128 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=15624 $Y=2940 $D=1
M295 91 87 129 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=15624 $Y=4884 $D=1
M296 Z<1> 90 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=16272 $Y=2940 $D=1
M297 Z<0> 91 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=16272 $Y=4884 $D=1
.ENDS
***************************************
