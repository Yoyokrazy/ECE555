#   Default technology Lef file
#   Created by correlating layers from PTF source [embedded corner "typical"] with SVRF rules "_rcxControl_calibre_asap7.rul_"

VERSION 5.7 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 2000 ;
END UNITS

LAYER Active
    TYPE ROUTING ;
    WIDTH 0.0118 ;
    PITCH 0.0388 ;
    DIRECTION VERTICAL ;
END Active

LAYER Activesd
    TYPE ROUTING ;
    WIDTH 0.0118 ;
    PITCH 0.0388 ;
    DIRECTION VERTICAL ;
END Activesd

LAYER Gate
    TYPE ROUTING ;
    WIDTH 0.021 ;
    PITCH 0.054 ;
    DIRECTION VERTICAL ;
END Gate

LAYER FGATE
    TYPE ROUTING ;
    WIDTH 0.021 ;
    PITCH 0.054 ;
    DIRECTION VERTICAL ;
END FGATE

LAYER SDT
    TYPE ROUTING ;
    WIDTH 0.0118 ;
    PITCH 0.054 ;
    DIRECTION VERTICAL ;
END SDT

LAYER LIG
    TYPE ROUTING ;
    WIDTH 0.016 ;
    PITCH 0.032 ;
    DIRECTION VERTICAL ;
END LIG

LAYER LISD
    TYPE ROUTING ;
    WIDTH 0.0118 ;
    PITCH 0.054 ;
    DIRECTION VERTICAL ;
END LISD

LAYER V0LISD
    TYPE CUT ;
END V0LISD

LAYER M1
    TYPE ROUTING ;
    WIDTH 0.018 ;
    PITCH 0.036 ;
    DIRECTION VERTICAL ;
END M1

LAYER V1
    TYPE CUT ;
END V1

LAYER M2
    TYPE ROUTING ;
    WIDTH 0.018 ;
    PITCH 0.036 ;
    DIRECTION VERTICAL ;
END M2

LAYER V2
    TYPE CUT ;
END V2

LAYER M3
    TYPE ROUTING ;
    WIDTH 0.018 ;
    PITCH 0.036 ;
    DIRECTION VERTICAL ;
END M3

LAYER V3
    TYPE CUT ;
END V3

LAYER M4
    TYPE ROUTING ;
    WIDTH 0.024 ;
    PITCH 0.048 ;
    DIRECTION VERTICAL ;
END M4

LAYER V4
    TYPE CUT ;
END V4

LAYER M5
    TYPE ROUTING ;
    WIDTH 0.024 ;
    PITCH 0.048 ;
    DIRECTION VERTICAL ;
END M5

LAYER V5
    TYPE CUT ;
END V5

LAYER M6
    TYPE ROUTING ;
    WIDTH 0.032 ;
    PITCH 0.064 ;
    DIRECTION VERTICAL ;
END M6

LAYER V6
    TYPE CUT ;
END V6

LAYER M7
    TYPE ROUTING ;
    WIDTH 0.032 ;
    PITCH 0.064 ;
    DIRECTION VERTICAL ;
END M7

LAYER V7
    TYPE CUT ;
END V7

LAYER M8
    TYPE ROUTING ;
    WIDTH 0.04 ;
    PITCH 0.08 ;
    DIRECTION VERTICAL ;
END M8

LAYER V8
    TYPE CUT ;
END V8

LAYER M9
    TYPE ROUTING ;
    WIDTH 0.04 ;
    PITCH 0.08 ;
    DIRECTION VERTICAL ;
END M9


#   Extra vias---

#   Via for layers FGATE and LIG
LAYER fvia_FGATE_LIG
    TYPE CUT ;
END fvia_FGATE_LIG

#   Via for layers LIG and M1
LAYER V0LIG
    TYPE CUT ;
END V0LIG

#   Via for layers SDT and LISD
LAYER COSD
    TYPE CUT ;
END COSD

#   Via for layers Gate and LIG
LAYER COG
    TYPE CUT ;
END COG

#   Via for layers Activesd and SDT
LAYER DIFF2SDT
    TYPE CUT ;
END DIFF2SDT

END LIBRARY
