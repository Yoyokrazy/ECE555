* SPICE NETLIST
***************************************

.SUBCKT NEURON VSS VDD X_1<0> X_0<0> W1_0<0> W1_0<1> W0_0<0> W0_0<1> X_1<1> X_0<1> CIN_0 W2_0<0> W2_0<1> W2_0<2> CIN_1 Z<2> Z<0> Z<1> COUT
** N=430 EP=19 IP=0 FDC=298
M0 11 X_1<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=972 $D=0
M1 VDD 4 15 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=1512 $D=0
M2 12 X_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=3456 $D=0
M3 VDD 6 16 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=3996 $D=0
M4 VDD W1_0<0> 11 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=972 $D=0
M5 142 W1_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=1512 $D=0
M6 VDD W0_0<0> 12 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=3456 $D=0
M7 143 W0_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=3996 $D=0
M8 15 X_1<1> 142 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=1512 $D=0
M9 16 X_0<1> 143 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=3996 $D=0
M10 19 11 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=756 $D=0
M11 20 12 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=3240 $D=0
M12 4 X_1<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=1512 $D=0
M13 6 X_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=3996 $D=0
M14 VDD W1_0<1> 4 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=1512 $D=0
M15 VDD W0_0<1> 6 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=3996 $D=0
M16 17 15 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=1512 $D=0
M17 18 16 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=3996 $D=0
M18 21 17 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=972 $D=0
M19 VDD 15 17 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=1512 $D=0
M20 22 18 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=3456 $D=0
M21 VDD 16 18 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=3996 $D=0
M22 VDD 19 21 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=972 $D=0
M23 VDD 20 22 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=3456 $D=0
M24 24 21 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=756 $D=0
M25 26 22 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=3240 $D=0
M26 29 20 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=972 $D=0
M27 VDD 23 34 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=1512 $D=0
M28 30 24 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=3456 $D=0
M29 VDD 25 35 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=3996 $D=0
M30 VDD 19 29 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=972 $D=0
M31 144 20 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=1512 $D=0
M32 VDD 26 30 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=3456 $D=0
M33 145 24 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=3996 $D=0
M34 34 19 144 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=1512 $D=0
M35 35 26 145 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=3996 $D=0
M36 VDD 27 Z<0> VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=5940 $D=0
M37 VDD 28 Z<1> VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=6588 $D=0
M38 47 29 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=756 $D=0
M39 48 30 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=3240 $D=0
M40 23 19 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=1512 $D=0
M41 25 26 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=3996 $D=0
M42 27 31 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=6156 $D=0
M43 28 32 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=6588 $D=0
M44 VDD 20 23 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=1512 $D=0
M45 VDD 24 25 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=3996 $D=0
M46 VDD 33 27 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=6156 $D=0
M47 VDD 31 28 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=6588 $D=0
M48 36 34 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=1512 $D=0
M49 37 35 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=3996 $D=0
M50 43 36 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5616 $Y=972 $D=0
M51 VDD 34 36 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=1512 $D=0
M52 44 37 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5616 $Y=3456 $D=0
M53 VDD 35 37 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=3996 $D=0
M54 VDD CIN_0 43 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5832 $Y=972 $D=0
M55 VDD 39 44 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5832 $Y=3456 $D=0
M56 VDD 40 31 VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=5940 $D=0
M57 VDD VDD Z<2> VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=6588 $D=0
M58 VDD 41 49 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=1512 $D=0
M59 VDD 42 50 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=3996 $D=0
M60 45 43 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=756 $D=0
M61 146 CIN_0 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=1512 $D=0
M62 46 44 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=3240 $D=0
M63 147 39 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=3996 $D=0
M64 49 36 146 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=1512 $D=0
M65 50 37 147 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=3996 $D=0
M66 119 45 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7128 $Y=972 $D=0
M67 120 46 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7128 $Y=3456 $D=0
M68 51 47 119 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=972 $D=0
M69 41 36 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=1512 $D=0
M70 52 48 120 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=3456 $D=0
M71 42 37 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=3996 $D=0
M72 VDD CIN_0 41 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7560 $Y=1512 $D=0
M73 VDD 39 42 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7560 $Y=3996 $D=0
M74 59 49 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=1512 $D=0
M75 60 50 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=3996 $D=0
M76 39 51 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7992 $Y=972 $D=0
M77 VDD 49 59 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=1512 $D=0
M78 61 52 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7992 $Y=3456 $D=0
M79 VDD 50 60 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=3996 $D=0
M80 62 W2_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=972 $D=0
M81 VDD 54 65 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=1512 $D=0
M82 63 W2_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=3456 $D=0
M83 VDD 56 66 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=3996 $D=0
M84 64 W2_0<2> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=5940 $D=0
M85 VDD 58 67 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=6480 $D=0
M86 VDD 59 62 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=972 $D=0
M87 148 W2_0<0> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=1512 $D=0
M88 VDD 60 63 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=3456 $D=0
M89 149 W2_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=3996 $D=0
M90 VDD 61 64 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=5940 $D=0
M91 150 W2_0<2> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=6480 $D=0
M92 65 59 148 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=1512 $D=0
M93 66 60 149 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=3996 $D=0
M94 67 61 150 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=6480 $D=0
M95 83 62 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=756 $D=0
M96 84 63 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=3240 $D=0
M97 85 64 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=5724 $D=0
M98 54 59 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=1512 $D=0
M99 56 60 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=3996 $D=0
M100 58 61 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=6480 $D=0
M101 VDD W2_0<0> 54 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=1512 $D=0
M102 VDD W2_0<1> 56 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=3996 $D=0
M103 VDD W2_0<2> 58 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=6480 $D=0
M104 68 65 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=1512 $D=0
M105 69 66 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=3996 $D=0
M106 70 67 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=6480 $D=0
M107 77 68 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=972 $D=0
M108 VDD 65 68 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=1512 $D=0
M109 78 69 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=3456 $D=0
M110 VDD 66 69 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=3996 $D=0
M111 79 70 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=5940 $D=0
M112 VDD 67 70 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=6480 $D=0
M113 VDD CIN_1 77 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=972 $D=0
M114 VDD 72 78 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=3456 $D=0
M115 VDD 73 79 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=5940 $D=0
M116 VDD 74 86 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=1512 $D=0
M117 VDD 75 87 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=3996 $D=0
M118 VDD 76 88 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=6480 $D=0
M119 80 77 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=756 $D=0
M120 151 CIN_1 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=1512 $D=0
M121 81 78 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=3240 $D=0
M122 152 72 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=3996 $D=0
M123 82 79 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=5724 $D=0
M124 153 73 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=6480 $D=0
M125 86 68 151 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=1512 $D=0
M126 87 69 152 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=3996 $D=0
M127 88 70 153 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=6480 $D=0
M128 127 80 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=972 $D=0
M129 128 81 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=3456 $D=0
M130 129 82 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=5940 $D=0
M131 89 83 127 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=972 $D=0
M132 74 68 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=1512 $D=0
M133 90 84 128 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=3456 $D=0
M134 75 69 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=3996 $D=0
M135 91 85 129 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=5940 $D=0
M136 76 70 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=6480 $D=0
M137 VDD CIN_1 74 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=1512 $D=0
M138 VDD 72 75 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=3996 $D=0
M139 VDD 73 76 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=6480 $D=0
M140 32 86 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=1512 $D=0
M141 33 87 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=3996 $D=0
M142 40 88 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=6480 $D=0
M143 72 89 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=972 $D=0
M144 VDD 86 32 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=1512 $D=0
M145 73 90 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=3456 $D=0
M146 VDD 87 33 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=3996 $D=0
M147 COUT 91 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=5940 $D=0
M148 VDD 88 40 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=6480 $D=0
M149 109 X_1<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=108 $D=1
M150 92 4 15 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=2052 $D=1
M151 110 X_0<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=2592 $D=1
M152 93 6 16 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=4536 $D=1
M153 11 W1_0<0> 109 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=108 $D=1
M154 VSS W1_0<1> 92 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=2052 $D=1
M155 12 W0_0<0> 110 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=2592 $D=1
M156 VSS W0_0<1> 93 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=4536 $D=1
M157 92 X_1<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=2052 $D=1
M158 93 X_0<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=4536 $D=1
M159 19 11 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=108 $D=1
M160 20 12 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=2592 $D=1
M161 130 X_1<1> 4 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=2052 $D=1
M162 131 X_0<1> 6 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=4536 $D=1
M163 VSS W1_0<1> 130 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=2052 $D=1
M164 VSS W0_0<1> 131 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=4536 $D=1
M165 17 15 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=2052 $D=1
M166 18 16 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=4536 $D=1
M167 111 17 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=108 $D=1
M168 VSS 15 17 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=2052 $D=1
M169 112 18 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=2592 $D=1
M170 VSS 16 18 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=4536 $D=1
M171 21 19 111 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=108 $D=1
M172 22 20 112 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=2592 $D=1
M173 24 21 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=108 $D=1
M174 26 22 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=2592 $D=1
M175 113 20 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=108 $D=1
M176 95 23 34 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=2052 $D=1
M177 114 24 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=2592 $D=1
M178 96 25 35 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=4536 $D=1
M179 29 19 113 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4104 $Y=108 $D=1
M180 VSS 20 95 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=2052 $D=1
M181 30 26 114 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4104 $Y=2592 $D=1
M182 VSS 24 96 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=4536 $D=1
M183 95 19 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=2052 $D=1
M184 96 26 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=4536 $D=1
M185 VSS 27 Z<0> VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=5292 $D=1
M186 VSS 28 Z<1> VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=7236 $D=1
M187 47 29 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=108 $D=1
M188 48 30 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=2592 $D=1
M189 132 19 23 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4968 $Y=2052 $D=1
M190 133 26 25 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4968 $Y=4536 $D=1
M191 115 31 27 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4968 $Y=5292 $D=1
M192 116 32 28 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4968 $Y=7236 $D=1
M193 VSS 20 132 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5184 $Y=2052 $D=1
M194 VSS 24 133 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5184 $Y=4536 $D=1
M195 VSS 33 115 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5184 $Y=5292 $D=1
M196 VSS 31 116 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5184 $Y=7236 $D=1
M197 36 34 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=2052 $D=1
M198 37 35 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=4536 $D=1
M199 117 36 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5616 $Y=108 $D=1
M200 VSS 34 36 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=2052 $D=1
M201 118 37 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5616 $Y=2592 $D=1
M202 VSS 35 37 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=4536 $D=1
M203 43 CIN_0 117 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5832 $Y=108 $D=1
M204 44 39 118 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5832 $Y=2592 $D=1
M205 VSS 40 31 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=5292 $D=1
M206 VSS VDD Z<2> VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=7236 $D=1
M207 99 41 49 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=2052 $D=1
M208 100 42 50 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=4536 $D=1
M209 45 43 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=108 $D=1
M210 VSS CIN_0 99 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=2052 $D=1
M211 46 44 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=2592 $D=1
M212 VSS 39 100 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=4536 $D=1
M213 99 36 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=2052 $D=1
M214 100 37 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=4536 $D=1
M215 51 45 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7128 $Y=108 $D=1
M216 52 46 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7128 $Y=2592 $D=1
M217 VSS 47 51 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7344 $Y=108 $D=1
M218 134 36 41 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7344 $Y=2052 $D=1
M219 VSS 48 52 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7344 $Y=2592 $D=1
M220 135 37 42 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7344 $Y=4536 $D=1
M221 VSS CIN_0 134 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7560 $Y=2052 $D=1
M222 VSS 39 135 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7560 $Y=4536 $D=1
M223 59 49 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=2052 $D=1
M224 60 50 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=4536 $D=1
M225 39 51 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7992 $Y=108 $D=1
M226 VSS 49 59 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=2052 $D=1
M227 61 52 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7992 $Y=2592 $D=1
M228 VSS 50 60 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=4536 $D=1
M229 121 W2_0<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=108 $D=1
M230 102 54 65 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=2052 $D=1
M231 122 W2_0<1> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=2592 $D=1
M232 103 56 66 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=4536 $D=1
M233 123 W2_0<2> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=5076 $D=1
M234 104 58 67 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=7020 $D=1
M235 62 59 121 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=108 $D=1
M236 VSS W2_0<0> 102 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=2052 $D=1
M237 63 60 122 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=2592 $D=1
M238 VSS W2_0<1> 103 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=4536 $D=1
M239 64 61 123 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=5076 $D=1
M240 VSS W2_0<2> 104 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=7020 $D=1
M241 102 59 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=2052 $D=1
M242 103 60 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=4536 $D=1
M243 104 61 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=7020 $D=1
M244 83 62 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=108 $D=1
M245 84 63 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=2592 $D=1
M246 85 64 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=5076 $D=1
M247 136 59 54 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=2052 $D=1
M248 137 60 56 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=4536 $D=1
M249 138 61 58 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=7020 $D=1
M250 VSS W2_0<0> 136 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=2052 $D=1
M251 VSS W2_0<1> 137 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=4536 $D=1
M252 VSS W2_0<2> 138 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=7020 $D=1
M253 68 65 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=2052 $D=1
M254 69 66 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=4536 $D=1
M255 70 67 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=7020 $D=1
M256 124 68 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=108 $D=1
M257 VSS 65 68 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=2052 $D=1
M258 125 69 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=2592 $D=1
M259 VSS 66 69 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=4536 $D=1
M260 126 70 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=5076 $D=1
M261 VSS 67 70 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=7020 $D=1
M262 77 CIN_1 124 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=108 $D=1
M263 78 72 125 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=2592 $D=1
M264 79 73 126 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=5076 $D=1
M265 105 74 86 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=2052 $D=1
M266 106 75 87 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=4536 $D=1
M267 107 76 88 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=7020 $D=1
M268 80 77 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=108 $D=1
M269 VSS CIN_1 105 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=2052 $D=1
M270 81 78 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=2592 $D=1
M271 VSS 72 106 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=4536 $D=1
M272 82 79 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=5076 $D=1
M273 VSS 73 107 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=7020 $D=1
M274 105 68 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=2052 $D=1
M275 106 69 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=4536 $D=1
M276 107 70 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=7020 $D=1
M277 89 80 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=108 $D=1
M278 90 81 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=2592 $D=1
M279 91 82 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=5076 $D=1
M280 VSS 83 89 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=108 $D=1
M281 139 68 74 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=2052 $D=1
M282 VSS 84 90 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=2592 $D=1
M283 140 69 75 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=4536 $D=1
M284 VSS 85 91 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=5076 $D=1
M285 141 70 76 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=7020 $D=1
M286 VSS CIN_1 139 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=2052 $D=1
M287 VSS 72 140 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=4536 $D=1
M288 VSS 73 141 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=7020 $D=1
M289 32 86 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=2052 $D=1
M290 33 87 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=4536 $D=1
M291 40 88 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=7020 $D=1
M292 72 89 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=108 $D=1
M293 VSS 86 32 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=2052 $D=1
M294 73 90 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=2592 $D=1
M295 VSS 87 33 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=4536 $D=1
M296 COUT 91 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=5076 $D=1
M297 VSS 88 40 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=7020 $D=1
.ENDS
***************************************
