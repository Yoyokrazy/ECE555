* SPICE NETLIST
***************************************

.SUBCKT NEURON VSS VDD X_1<0> X_0<0> W1_0<0> W1_0<1> W0_0<0> W0_0<1> X_1<1> X_0<1> CIN_0 W2_0<0> W2_0<1> W2_0<2> CIN_1 Z<2> Z<0> Z<1> COUT
** N=430 EP=19 IP=0 FDC=298
M0 109 X_1<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=108 $D=1
M1 92 4 15 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=2052 $D=1
M2 110 X_0<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=2592 $D=1
M3 93 6 16 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=4536 $D=1
M4 11 W1_0<0> 109 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=108 $D=1
M5 VSS W1_0<1> 92 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=2052 $D=1
M6 12 W0_0<0> 110 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=2592 $D=1
M7 VSS W0_0<1> 93 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=4536 $D=1
M8 92 X_1<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=2052 $D=1
M9 93 X_0<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=4536 $D=1
M10 19 11 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=108 $D=1
M11 20 12 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=2592 $D=1
M12 130 X_1<1> 4 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=2052 $D=1
M13 131 X_0<1> 6 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=4536 $D=1
M14 VSS W1_0<1> 130 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=2052 $D=1
M15 VSS W0_0<1> 131 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=4536 $D=1
M16 17 15 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=2052 $D=1
M17 18 16 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=4536 $D=1
M18 111 17 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=108 $D=1
M19 VSS 15 17 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=2052 $D=1
M20 112 18 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=2592 $D=1
M21 VSS 16 18 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=4536 $D=1
M22 21 19 111 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=108 $D=1
M23 22 20 112 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=2592 $D=1
M24 24 21 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=108 $D=1
M25 26 22 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=2592 $D=1
M26 113 20 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=108 $D=1
M27 95 23 34 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=2052 $D=1
M28 114 24 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=2592 $D=1
M29 96 25 35 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=4536 $D=1
M30 29 19 113 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4104 $Y=108 $D=1
M31 VSS 20 95 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=2052 $D=1
M32 30 26 114 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4104 $Y=2592 $D=1
M33 VSS 24 96 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=4536 $D=1
M34 95 19 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=2052 $D=1
M35 96 26 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=4536 $D=1
M36 VSS 27 Z<0> VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=5292 $D=1
M37 VSS 28 Z<1> VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=7236 $D=1
M38 47 29 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=108 $D=1
M39 48 30 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=2592 $D=1
M40 132 19 23 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4968 $Y=2052 $D=1
M41 133 26 25 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4968 $Y=4536 $D=1
M42 115 31 27 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4968 $Y=5292 $D=1
M43 116 32 28 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4968 $Y=7236 $D=1
M44 VSS 20 132 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5184 $Y=2052 $D=1
M45 VSS 24 133 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5184 $Y=4536 $D=1
M46 VSS 33 115 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5184 $Y=5292 $D=1
M47 VSS 31 116 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5184 $Y=7236 $D=1
M48 36 34 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=2052 $D=1
M49 37 35 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=4536 $D=1
M50 117 36 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5616 $Y=108 $D=1
M51 VSS 34 36 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=2052 $D=1
M52 118 37 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5616 $Y=2592 $D=1
M53 VSS 35 37 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=4536 $D=1
M54 43 CIN_0 117 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5832 $Y=108 $D=1
M55 44 39 118 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=5832 $Y=2592 $D=1
M56 VSS 40 31 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=5292 $D=1
M57 VSS VDD Z<2> VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=7236 $D=1
M58 99 41 49 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=2052 $D=1
M59 100 42 50 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=4536 $D=1
M60 45 43 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=108 $D=1
M61 VSS CIN_0 99 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=2052 $D=1
M62 46 44 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=2592 $D=1
M63 VSS 39 100 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=4536 $D=1
M64 99 36 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=2052 $D=1
M65 100 37 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=4536 $D=1
M66 51 45 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7128 $Y=108 $D=1
M67 52 46 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7128 $Y=2592 $D=1
M68 VSS 47 51 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7344 $Y=108 $D=1
M69 134 36 41 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7344 $Y=2052 $D=1
M70 VSS 48 52 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7344 $Y=2592 $D=1
M71 135 37 42 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7344 $Y=4536 $D=1
M72 VSS CIN_0 134 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7560 $Y=2052 $D=1
M73 VSS 39 135 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7560 $Y=4536 $D=1
M74 59 49 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=2052 $D=1
M75 60 50 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=4536 $D=1
M76 39 51 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7992 $Y=108 $D=1
M77 VSS 49 59 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=2052 $D=1
M78 61 52 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=7992 $Y=2592 $D=1
M79 VSS 50 60 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=4536 $D=1
M80 121 W2_0<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=108 $D=1
M81 102 54 65 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=2052 $D=1
M82 122 W2_0<1> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=2592 $D=1
M83 103 56 66 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=4536 $D=1
M84 123 W2_0<2> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9152 $Y=5076 $D=1
M85 104 58 67 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=7020 $D=1
M86 62 59 121 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=108 $D=1
M87 VSS W2_0<0> 102 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=2052 $D=1
M88 63 60 122 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=2592 $D=1
M89 VSS W2_0<1> 103 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=4536 $D=1
M90 64 61 123 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=9368 $Y=5076 $D=1
M91 VSS W2_0<2> 104 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=7020 $D=1
M92 102 59 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=2052 $D=1
M93 103 60 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=4536 $D=1
M94 104 61 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=7020 $D=1
M95 83 62 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=108 $D=1
M96 84 63 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=2592 $D=1
M97 85 64 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=5076 $D=1
M98 136 59 54 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=2052 $D=1
M99 137 60 56 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=4536 $D=1
M100 138 61 58 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10232 $Y=7020 $D=1
M101 VSS W2_0<0> 136 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=2052 $D=1
M102 VSS W2_0<1> 137 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=4536 $D=1
M103 VSS W2_0<2> 138 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10448 $Y=7020 $D=1
M104 68 65 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=2052 $D=1
M105 69 66 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=4536 $D=1
M106 70 67 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=7020 $D=1
M107 124 68 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=108 $D=1
M108 VSS 65 68 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=2052 $D=1
M109 125 69 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=2592 $D=1
M110 VSS 66 69 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=4536 $D=1
M111 126 70 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10880 $Y=5076 $D=1
M112 VSS 67 70 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=7020 $D=1
M113 77 CIN_1 124 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=108 $D=1
M114 78 72 125 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=2592 $D=1
M115 79 73 126 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11096 $Y=5076 $D=1
M116 105 74 86 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=2052 $D=1
M117 106 75 87 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=4536 $D=1
M118 107 76 88 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=7020 $D=1
M119 80 77 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=108 $D=1
M120 VSS CIN_1 105 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=2052 $D=1
M121 81 78 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=2592 $D=1
M122 VSS 72 106 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=4536 $D=1
M123 82 79 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=5076 $D=1
M124 VSS 73 107 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=7020 $D=1
M125 105 68 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=2052 $D=1
M126 106 69 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=4536 $D=1
M127 107 70 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=7020 $D=1
M128 89 80 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=108 $D=1
M129 90 81 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=2592 $D=1
M130 91 82 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12392 $Y=5076 $D=1
M131 VSS 83 89 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=108 $D=1
M132 139 68 74 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=2052 $D=1
M133 VSS 84 90 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=2592 $D=1
M134 140 69 75 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=4536 $D=1
M135 VSS 85 91 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=12608 $Y=5076 $D=1
M136 141 70 76 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12608 $Y=7020 $D=1
M137 VSS CIN_1 139 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=2052 $D=1
M138 VSS 72 140 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=4536 $D=1
M139 VSS 73 141 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=12824 $Y=7020 $D=1
M140 32 86 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=2052 $D=1
M141 33 87 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=4536 $D=1
M142 40 88 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=7020 $D=1
M143 72 89 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=108 $D=1
M144 VSS 86 32 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=2052 $D=1
M145 73 90 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=2592 $D=1
M146 VSS 87 33 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=4536 $D=1
M147 COUT 91 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=13256 $Y=5076 $D=1
M148 VSS 88 40 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=7020 $D=1
M149 11 X_1<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=972 $D=0
M150 VDD 4 15 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=1512 $D=0
M151 12 X_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=3456 $D=0
M152 VDD 6 16 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=3996 $D=0
M153 VDD W1_0<0> 11 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=972 $D=0
M154 142 W1_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=1512 $D=0
M155 VDD W0_0<0> 12 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=3456 $D=0
M156 143 W0_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=3996 $D=0
M157 15 X_1<1> 142 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=1512 $D=0
M158 16 X_0<1> 143 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=3996 $D=0
M159 19 11 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=756 $D=0
M160 20 12 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=3240 $D=0
M161 4 X_1<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=1512 $D=0
M162 6 X_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=3996 $D=0
M163 VDD W1_0<1> 4 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=1512 $D=0
M164 VDD W0_0<1> 6 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=3996 $D=0
M165 17 15 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=1512 $D=0
M166 18 16 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=3996 $D=0
M167 21 17 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=972 $D=0
M168 VDD 15 17 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=1512 $D=0
M169 22 18 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=3456 $D=0
M170 VDD 16 18 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=3996 $D=0
M171 VDD 19 21 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=972 $D=0
M172 VDD 20 22 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=3456 $D=0
M173 24 21 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=756 $D=0
M174 26 22 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=3240 $D=0
M175 29 20 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=972 $D=0
M176 VDD 23 34 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=1512 $D=0
M177 30 24 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=3456 $D=0
M178 VDD 25 35 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=3996 $D=0
M179 VDD 19 29 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=972 $D=0
M180 144 20 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=1512 $D=0
M181 VDD 26 30 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=3456 $D=0
M182 145 24 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=3996 $D=0
M183 34 19 144 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=1512 $D=0
M184 35 26 145 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=3996 $D=0
M185 VDD 27 Z<0> VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=5940 $D=0
M186 VDD 28 Z<1> VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4320 $Y=6588 $D=0
M187 47 29 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=756 $D=0
M188 48 30 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4752 $Y=3240 $D=0
M189 23 19 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=1512 $D=0
M190 25 26 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=3996 $D=0
M191 27 31 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=6156 $D=0
M192 28 32 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4968 $Y=6588 $D=0
M193 VDD 20 23 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=1512 $D=0
M194 VDD 24 25 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=3996 $D=0
M195 VDD 33 27 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=6156 $D=0
M196 VDD 31 28 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5184 $Y=6588 $D=0
M197 36 34 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=1512 $D=0
M198 37 35 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5400 $Y=3996 $D=0
M199 43 36 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5616 $Y=972 $D=0
M200 VDD 34 36 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=1512 $D=0
M201 44 37 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5616 $Y=3456 $D=0
M202 VDD 35 37 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5616 $Y=3996 $D=0
M203 VDD CIN_0 43 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5832 $Y=972 $D=0
M204 VDD 39 44 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5832 $Y=3456 $D=0
M205 VDD 40 31 VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=5940 $D=0
M206 VDD VDD Z<2> VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6128 $Y=6588 $D=0
M207 VDD 41 49 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=1512 $D=0
M208 VDD 42 50 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6264 $Y=3996 $D=0
M209 45 43 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=756 $D=0
M210 146 CIN_0 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=1512 $D=0
M211 46 44 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=6480 $Y=3240 $D=0
M212 147 39 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6480 $Y=3996 $D=0
M213 49 36 146 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=1512 $D=0
M214 50 37 147 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6696 $Y=3996 $D=0
M215 119 45 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7128 $Y=972 $D=0
M216 120 46 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7128 $Y=3456 $D=0
M217 51 47 119 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=972 $D=0
M218 41 36 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=1512 $D=0
M219 52 48 120 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=3456 $D=0
M220 42 37 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7344 $Y=3996 $D=0
M221 VDD CIN_0 41 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7560 $Y=1512 $D=0
M222 VDD 39 42 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7560 $Y=3996 $D=0
M223 59 49 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=1512 $D=0
M224 60 50 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7776 $Y=3996 $D=0
M225 39 51 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7992 $Y=972 $D=0
M226 VDD 49 59 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=1512 $D=0
M227 61 52 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7992 $Y=3456 $D=0
M228 VDD 50 60 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7992 $Y=3996 $D=0
M229 62 W2_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=972 $D=0
M230 VDD 54 65 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=1512 $D=0
M231 63 W2_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=3456 $D=0
M232 VDD 56 66 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=3996 $D=0
M233 64 W2_0<2> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9152 $Y=5940 $D=0
M234 VDD 58 67 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9152 $Y=6480 $D=0
M235 VDD 59 62 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=972 $D=0
M236 148 W2_0<0> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=1512 $D=0
M237 VDD 60 63 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=3456 $D=0
M238 149 W2_0<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=3996 $D=0
M239 VDD 61 64 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=9368 $Y=5940 $D=0
M240 150 W2_0<2> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9368 $Y=6480 $D=0
M241 65 59 148 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=1512 $D=0
M242 66 60 149 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=3996 $D=0
M243 67 61 150 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=9584 $Y=6480 $D=0
M244 83 62 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=756 $D=0
M245 84 63 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=3240 $D=0
M246 85 64 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=10016 $Y=5724 $D=0
M247 54 59 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=1512 $D=0
M248 56 60 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=3996 $D=0
M249 58 61 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10232 $Y=6480 $D=0
M250 VDD W2_0<0> 54 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=1512 $D=0
M251 VDD W2_0<1> 56 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=3996 $D=0
M252 VDD W2_0<2> 58 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10448 $Y=6480 $D=0
M253 68 65 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=1512 $D=0
M254 69 66 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=3996 $D=0
M255 70 67 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10664 $Y=6480 $D=0
M256 77 68 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=972 $D=0
M257 VDD 65 68 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=1512 $D=0
M258 78 69 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=3456 $D=0
M259 VDD 66 69 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=3996 $D=0
M260 79 70 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=10880 $Y=5940 $D=0
M261 VDD 67 70 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=10880 $Y=6480 $D=0
M262 VDD CIN_1 77 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=972 $D=0
M263 VDD 72 78 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=3456 $D=0
M264 VDD 73 79 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=11096 $Y=5940 $D=0
M265 VDD 74 86 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=1512 $D=0
M266 VDD 75 87 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=3996 $D=0
M267 VDD 76 88 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11528 $Y=6480 $D=0
M268 80 77 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=756 $D=0
M269 151 CIN_1 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=1512 $D=0
M270 81 78 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=3240 $D=0
M271 152 72 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=3996 $D=0
M272 82 79 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=11744 $Y=5724 $D=0
M273 153 73 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11744 $Y=6480 $D=0
M274 86 68 151 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=1512 $D=0
M275 87 69 152 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=3996 $D=0
M276 88 70 153 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=11960 $Y=6480 $D=0
M277 127 80 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=972 $D=0
M278 128 81 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=3456 $D=0
M279 129 82 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12392 $Y=5940 $D=0
M280 89 83 127 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=972 $D=0
M281 74 68 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=1512 $D=0
M282 90 84 128 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=3456 $D=0
M283 75 69 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=3996 $D=0
M284 91 85 129 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=5940 $D=0
M285 76 70 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12608 $Y=6480 $D=0
M286 VDD CIN_1 74 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=1512 $D=0
M287 VDD 72 75 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=3996 $D=0
M288 VDD 73 76 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=12824 $Y=6480 $D=0
M289 32 86 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=1512 $D=0
M290 33 87 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=3996 $D=0
M291 40 88 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13040 $Y=6480 $D=0
M292 72 89 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=972 $D=0
M293 VDD 86 32 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=1512 $D=0
M294 73 90 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=3456 $D=0
M295 VDD 87 33 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=3996 $D=0
M296 COUT 91 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=13256 $Y=5940 $D=0
M297 VDD 88 40 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=13256 $Y=6480 $D=0
.ENDS
***************************************
