* SPICE NETLIST
***************************************

.SUBCKT ADD3 VSS VDD IN_1<0> IN_1<1> IN_1<2> IN_0<0> IN_0<1> IN_0<2> CIN SUM<0> SUM<1> SUM<2> COUT
** N=190 EP=13 IP=0 FDC=138
M0 53 IN_1<0> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=104 $D=1
M1 43 4 15 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=2048 $D=1
M2 54 IN_1<1> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=2588 $D=1
M3 44 6 16 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=4532 $D=1
M4 55 IN_1<2> VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=432 $Y=5072 $D=1
M5 45 8 17 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=7016 $D=1
M6 12 IN_0<0> 53 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=104 $D=1
M7 VSS IN_1<0> 43 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=2048 $D=1
M8 13 IN_0<1> 54 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=2588 $D=1
M9 VSS IN_1<1> 44 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=4532 $D=1
M10 14 IN_0<2> 55 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=648 $Y=5072 $D=1
M11 VSS IN_1<2> 45 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=7016 $D=1
M12 43 IN_0<0> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=2048 $D=1
M13 44 IN_0<1> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=4532 $D=1
M14 45 IN_0<2> VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=7016 $D=1
M15 33 12 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=104 $D=1
M16 34 13 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=2588 $D=1
M17 35 14 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=5072 $D=1
M18 62 IN_0<0> 4 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=2048 $D=1
M19 63 IN_0<1> 6 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=4532 $D=1
M20 64 IN_0<2> 8 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1512 $Y=7016 $D=1
M21 VSS IN_1<0> 62 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=2048 $D=1
M22 VSS IN_1<1> 63 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=4532 $D=1
M23 VSS IN_1<2> 64 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1728 $Y=7016 $D=1
M24 18 15 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=2048 $D=1
M25 19 16 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=4532 $D=1
M26 20 17 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=7016 $D=1
M27 56 18 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=104 $D=1
M28 VSS 15 18 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=2048 $D=1
M29 57 19 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=2588 $D=1
M30 VSS 16 19 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=4532 $D=1
M31 58 20 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2160 $Y=5072 $D=1
M32 VSS 17 20 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=7016 $D=1
M33 27 CIN 56 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=104 $D=1
M34 28 22 57 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=2588 $D=1
M35 29 23 58 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=2376 $Y=5072 $D=1
M36 46 24 36 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2808 $Y=2048 $D=1
M37 47 25 37 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2808 $Y=4532 $D=1
M38 48 26 38 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2808 $Y=7016 $D=1
M39 30 27 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=104 $D=1
M40 VSS CIN 46 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3024 $Y=2048 $D=1
M41 31 28 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=2588 $D=1
M42 VSS 22 47 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3024 $Y=4532 $D=1
M43 32 29 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=5072 $D=1
M44 VSS 23 48 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3024 $Y=7016 $D=1
M45 46 18 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3240 $Y=2048 $D=1
M46 47 19 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3240 $Y=4532 $D=1
M47 48 20 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3240 $Y=7016 $D=1
M48 39 30 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3672 $Y=104 $D=1
M49 40 31 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3672 $Y=2588 $D=1
M50 41 32 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3672 $Y=5072 $D=1
M51 VSS 33 39 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=104 $D=1
M52 65 18 24 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=2048 $D=1
M53 VSS 34 40 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=2588 $D=1
M54 66 19 25 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=4532 $D=1
M55 VSS 35 41 VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3888 $Y=5072 $D=1
M56 67 20 26 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3888 $Y=7016 $D=1
M57 VSS CIN 65 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=2048 $D=1
M58 VSS 22 66 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=4532 $D=1
M59 VSS 23 67 VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4104 $Y=7016 $D=1
M60 SUM<0> 36 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=2048 $D=1
M61 SUM<1> 37 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=4532 $D=1
M62 SUM<2> 38 VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=7016 $D=1
M63 22 39 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4536 $Y=104 $D=1
M64 VSS 36 SUM<0> VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4536 $Y=2048 $D=1
M65 23 40 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4536 $Y=2588 $D=1
M66 VSS 37 SUM<1> VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4536 $Y=4532 $D=1
M67 COUT 41 VSS VSS nmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=4536 $Y=5072 $D=1
M68 VSS 38 SUM<2> VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4536 $Y=7016 $D=1
M69 12 IN_1<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=968 $D=0
M70 VDD 4 15 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=1508 $D=0
M71 13 IN_1<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=3452 $D=0
M72 VDD 6 16 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=3992 $D=0
M73 14 IN_1<2> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=432 $Y=5936 $D=0
M74 VDD 8 17 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=432 $Y=6476 $D=0
M75 VDD IN_0<0> 12 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=968 $D=0
M76 68 IN_1<0> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=1508 $D=0
M77 VDD IN_0<1> 13 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=3452 $D=0
M78 69 IN_1<1> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=3992 $D=0
M79 VDD IN_0<2> 14 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=648 $Y=5936 $D=0
M80 70 IN_1<2> VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=648 $Y=6476 $D=0
M81 15 IN_0<0> 68 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=1508 $D=0
M82 16 IN_0<1> 69 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=3992 $D=0
M83 17 IN_0<2> 70 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=864 $Y=6476 $D=0
M84 33 12 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=752 $D=0
M85 34 13 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=3236 $D=0
M86 35 14 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=1296 $Y=5720 $D=0
M87 4 IN_0<0> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=1508 $D=0
M88 6 IN_0<1> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=3992 $D=0
M89 8 IN_0<2> VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1512 $Y=6476 $D=0
M90 VDD IN_1<0> 4 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=1508 $D=0
M91 VDD IN_1<1> 6 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=3992 $D=0
M92 VDD IN_1<2> 8 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1728 $Y=6476 $D=0
M93 18 15 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=1508 $D=0
M94 19 16 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=3992 $D=0
M95 20 17 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1944 $Y=6476 $D=0
M96 27 18 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=968 $D=0
M97 VDD 15 18 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=1508 $D=0
M98 28 19 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=3452 $D=0
M99 VDD 16 19 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=3992 $D=0
M100 29 20 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2160 $Y=5936 $D=0
M101 VDD 17 20 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2160 $Y=6476 $D=0
M102 VDD CIN 27 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=968 $D=0
M103 VDD 22 28 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=3452 $D=0
M104 VDD 23 29 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2376 $Y=5936 $D=0
M105 VDD 24 36 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2808 $Y=1508 $D=0
M106 VDD 25 37 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2808 $Y=3992 $D=0
M107 VDD 26 38 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2808 $Y=6476 $D=0
M108 30 27 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=752 $D=0
M109 71 CIN VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3024 $Y=1508 $D=0
M110 31 28 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=3236 $D=0
M111 72 22 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3024 $Y=3992 $D=0
M112 32 29 VDD VDD pmos_rvt L=2e-08 W=1.08e-07 nfin=4 $X=3024 $Y=5720 $D=0
M113 73 23 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3024 $Y=6476 $D=0
M114 36 18 71 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3240 $Y=1508 $D=0
M115 37 19 72 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3240 $Y=3992 $D=0
M116 38 20 73 VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3240 $Y=6476 $D=0
M117 59 30 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3672 $Y=968 $D=0
M118 60 31 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3672 $Y=3452 $D=0
M119 61 32 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3672 $Y=5936 $D=0
M120 39 33 59 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=968 $D=0
M121 24 18 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=1508 $D=0
M122 40 34 60 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=3452 $D=0
M123 25 19 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=3992 $D=0
M124 41 35 61 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=5936 $D=0
M125 26 20 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3888 $Y=6476 $D=0
M126 VDD CIN 24 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=1508 $D=0
M127 VDD 22 25 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=3992 $D=0
M128 VDD 23 26 VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4104 $Y=6476 $D=0
M129 SUM<0> 36 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=1508 $D=0
M130 SUM<1> 37 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=3992 $D=0
M131 SUM<2> 38 VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4320 $Y=6476 $D=0
M132 22 39 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4536 $Y=968 $D=0
M133 VDD 36 SUM<0> VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4536 $Y=1508 $D=0
M134 23 40 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4536 $Y=3452 $D=0
M135 VDD 37 SUM<1> VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4536 $Y=3992 $D=0
M136 COUT 41 VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4536 $Y=5936 $D=0
M137 VDD 38 SUM<2> VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4536 $Y=6476 $D=0
.ENDS
***************************************
